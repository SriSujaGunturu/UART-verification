package final_pkg;
   import uvm_pkg::*;   
 
   `include "uvm_macros.svh"
   `include "timescale.v"
   `include "transaction.sv"
   `include "source_cfg.sv"
   `include "env_config.sv"
   `include "base_sequence.sv"
   `include "driver.sv"
   `include "monitor.sv"
   `include "sequencer.sv"
   `include "agent.sv"
   `include "agent_top.sv"
   `include "scoreboard.sv"
   `include "virtual_seqr.sv"
   `include "virtual_seq.sv"
   `include "environment.sv"
   `include "base_test.sv"

endpackage
